library ieee;
use ieee.std_logic_1164.all;

entity Comparador_e is
	port(
			en	         : in std_logic;
			a				: in std_logic;
			b 				: in std_logic_vector(18 downto 0);
			ls				: out std_logic
		 );
end Comparador_e;

architecture arq1 of Comparador_e is
begin
	
end arq1;