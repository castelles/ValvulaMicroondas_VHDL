library ieee;
use ieee.std_logic_1164.all;

entity One_delay is
  port (
    d  : in  std_logic;
    q  : out std_logic;
    clk   : in  std_logic
  );
end One_delay;

architecture onedelay_arc of One_delay is
begin

end onedelay_arc;